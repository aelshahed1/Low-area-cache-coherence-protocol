//4-bit alu functions

`define FNONE 4'b0000
`define FADD 4'b0001 
`define FSUB 4'b0010
`define FMULT 4'b0011
`define FAND 4'b0100
`define FOR 4'b0101
`define FXOR 4'b0110
`define FSLL 4'b0111
`define FSRL 4'b1000
`define FSRA 4'b1001
`define FSLT 4'b1010
`define FSLTU 4'b1011
`define FMULTH 4'b1100 

